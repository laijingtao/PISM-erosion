netcdf paleo_modifier {
dimensions:
	time = 1 ;
	tbnds = 2 ;
variables:
	float time(time) ;
		time:long_name = "Time (years before present)" ;
		time:standard_name = "time" ;
		time:units = "years since 1-1-1" ;
		time:calendar = "365_day" ;
		time:bounds = "time_bnds" ;
	float time_bnds(time, tbnds) ;
	float frac_P(time) ;
	float delta_T(time) ;
		delta_T:units = "Kelvin" ;
data:

 frac_P = 1 ;
 delta_T = 0 ;

 time = 0 ;
 time_bnds = -1000000, 1000000 ;
}
